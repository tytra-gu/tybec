library verilog;
use verilog.vl_types.all;
entity krnl_vadd_rtl_int is
    generic(
        C_S_AXI_CONTROL_DATA_WIDTH: integer := 32;
        C_S_AXI_CONTROL_ADDR_WIDTH: integer := 6;
        C_M_AXI_GMEM_ID_WIDTH: integer := 1;
        C_M_AXI_GMEM_ADDR_WIDTH: integer := 64;
        C_M_AXI_GMEM_DATA_WIDTH: integer := 32
    );
    port(
        ap_clk          : in     vl_logic;
        ap_rst_n        : in     vl_logic;
        m_axi_gmem_AWVALID: out    vl_logic;
        m_axi_gmem_AWREADY: in     vl_logic;
        m_axi_gmem_AWADDR: out    vl_logic_vector;
        m_axi_gmem_AWID : out    vl_logic_vector;
        m_axi_gmem_AWLEN: out    vl_logic_vector(7 downto 0);
        m_axi_gmem_AWSIZE: out    vl_logic_vector(2 downto 0);
        m_axi_gmem_AWBURST: out    vl_logic_vector(1 downto 0);
        m_axi_gmem_AWLOCK: out    vl_logic_vector(1 downto 0);
        m_axi_gmem_AWCACHE: out    vl_logic_vector(3 downto 0);
        m_axi_gmem_AWPROT: out    vl_logic_vector(2 downto 0);
        m_axi_gmem_AWQOS: out    vl_logic_vector(3 downto 0);
        m_axi_gmem_AWREGION: out    vl_logic_vector(3 downto 0);
        m_axi_gmem_WVALID: out    vl_logic;
        m_axi_gmem_WREADY: in     vl_logic;
        m_axi_gmem_WDATA: out    vl_logic_vector;
        m_axi_gmem_WSTRB: out    vl_logic_vector;
        m_axi_gmem_WLAST: out    vl_logic;
        m_axi_gmem_ARVALID: out    vl_logic;
        m_axi_gmem_ARREADY: in     vl_logic;
        m_axi_gmem_ARADDR: out    vl_logic_vector;
        m_axi_gmem_ARID : out    vl_logic_vector;
        m_axi_gmem_ARLEN: out    vl_logic_vector(7 downto 0);
        m_axi_gmem_ARSIZE: out    vl_logic_vector(2 downto 0);
        m_axi_gmem_ARBURST: out    vl_logic_vector(1 downto 0);
        m_axi_gmem_ARLOCK: out    vl_logic_vector(1 downto 0);
        m_axi_gmem_ARCACHE: out    vl_logic_vector(3 downto 0);
        m_axi_gmem_ARPROT: out    vl_logic_vector(2 downto 0);
        m_axi_gmem_ARQOS: out    vl_logic_vector(3 downto 0);
        m_axi_gmem_ARREGION: out    vl_logic_vector(3 downto 0);
        m_axi_gmem_RVALID: in     vl_logic;
        m_axi_gmem_RREADY: out    vl_logic;
        m_axi_gmem_RDATA: in     vl_logic_vector;
        m_axi_gmem_RLAST: in     vl_logic;
        m_axi_gmem_RID  : in     vl_logic_vector;
        m_axi_gmem_RRESP: in     vl_logic_vector(1 downto 0);
        m_axi_gmem_BVALID: in     vl_logic;
        m_axi_gmem_BREADY: out    vl_logic;
        m_axi_gmem_BRESP: in     vl_logic_vector(1 downto 0);
        m_axi_gmem_BID  : in     vl_logic_vector;
        s_axi_control_AWVALID: in     vl_logic;
        s_axi_control_AWREADY: out    vl_logic;
        s_axi_control_AWADDR: in     vl_logic_vector;
        s_axi_control_WVALID: in     vl_logic;
        s_axi_control_WREADY: out    vl_logic;
        s_axi_control_WDATA: in     vl_logic_vector;
        s_axi_control_WSTRB: in     vl_logic_vector;
        s_axi_control_ARVALID: in     vl_logic;
        s_axi_control_ARREADY: out    vl_logic;
        s_axi_control_ARADDR: in     vl_logic_vector;
        s_axi_control_RVALID: out    vl_logic;
        s_axi_control_RREADY: in     vl_logic;
        s_axi_control_RDATA: out    vl_logic_vector;
        s_axi_control_RRESP: out    vl_logic_vector(1 downto 0);
        s_axi_control_BVALID: out    vl_logic;
        s_axi_control_BREADY: in     vl_logic;
        s_axi_control_BRESP: out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_S_AXI_CONTROL_DATA_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of C_S_AXI_CONTROL_ADDR_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of C_M_AXI_GMEM_ID_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of C_M_AXI_GMEM_ADDR_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of C_M_AXI_GMEM_DATA_WIDTH : constant is 2;
end krnl_vadd_rtl_int;
